module net_write_tracker(
    aclk,
    aresetn,
    
    
    
    
    );
    
    
endmodule
